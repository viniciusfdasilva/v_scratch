module mymodule

pub const golden_ratio = 1.61803

fn calc(){
	println(mymodule.golden_ratio)
}
