module sample

@[noinit]
pub struct Information{
	pub:
		data string
}

pub fn new_information(data string) !Information{

	if data.len == 0 || data.len > 100{
		return error('data must be between 1 and 100 characters')
	}else{
		return Information{
			data: data
		}
	}
}